LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY Main IS
GENERIC (N:integer:=16);
Port(
	clk,rst : IN std_logic
);
END Main;

ARCHITECTURE ArchMain OF Main IS
BEGIN

END ArchMain;